module riscv_core #(
) (
);
	
endmodule