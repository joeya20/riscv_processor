module control_unit (

);

	
endmodule : control_unit