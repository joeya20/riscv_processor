module riscv_top (
	input clk_i
);
	



endmodule