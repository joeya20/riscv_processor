//top level
module riscv_top (
	input clk_i
);
	
riscv_core core(

);

mem inst_mem(

);

mem data_mem(
	
);

endmodule